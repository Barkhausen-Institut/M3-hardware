
parameter MODID_TILE0  = 8'h04,
parameter MODID_TILE1  = 8'h05,
parameter MODID_TILE2  = 8'h06,
parameter MODID_TILE3  = 8'h24,
parameter MODID_TILE4  = 8'h25,
parameter MODID_TILE5  = 8'h26,
parameter MODID_TILE6  = 8'h00,
parameter MODID_TILE7  = 8'h01,
parameter MODID_TILE8  = 8'h02,
parameter MODID_TILE9  = 8'h20,
parameter MODID_TILE10 = 8'h21,
parameter MODID_TILE11 = 8'h22,

parameter MODID_PM0 = MODID_TILE2,
parameter MODID_PM1 = MODID_TILE4,
parameter MODID_PM2 = MODID_TILE5,
parameter MODID_PM3 = MODID_TILE6,
parameter MODID_PM4 = MODID_TILE7,
parameter MODID_PM5 = MODID_TILE8,
parameter MODID_PM6 = MODID_TILE9,
parameter MODID_PM7 = MODID_TILE10,

parameter MODID_UART  = MODID_TILE0,
parameter MODID_ETH   = MODID_TILE1,
parameter MODID_DRAM1 = MODID_TILE3,
parameter MODID_DRAM2 = MODID_TILE11,


parameter MODID_ROUTER0 = 8'h07,
parameter MODID_ROUTER1 = 8'h27,
parameter MODID_ROUTER2 = 8'h03,
parameter MODID_ROUTER3 = 8'h23
