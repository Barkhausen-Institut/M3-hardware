
//select PM type
//0: no PM
//1: Rocket
//2: Boom
//3: Ethernet FMC
parameter PM_TYPE_NONE     = 0,
parameter PM_TYPE_ROCKET   = 1,
parameter PM_TYPE_BOOM     = 2,
parameter PM_TYPE_ETHFMC   = 3,
parameter PM_TYPE_ACC      = 4
