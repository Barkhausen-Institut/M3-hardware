
parameter DDR4_STATUS_SIZE = 3,

parameter DDR4_ADDR_SHIFT = 6,

parameter DDR4_APP_CMD_WIDTH = 3,
parameter DDR4_APP_ADDR_WIDTH = 28,
parameter DDR4_APP_DATA_WIDTH = 640,
parameter DDR4_APP_DATA_CUT_WIDTH = 512
