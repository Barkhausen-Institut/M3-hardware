
parameter CHIPID_HOST  = {NOC_CHIPID_SIZE{1'b1}}

